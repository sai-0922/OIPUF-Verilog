`include "MUX2to1_group.v"

module lines4_stages64_diff(  
(* DONT_TOUCH= "TRUE" *)input itriger,     
(* DONT_TOUCH= "TRUE" *)input  [63 :0] iC, //   No. of challenge bits i.e., n stages
(* DONT_TOUCH= "TRUE" *)output [3 :0] oTP //    No. of output bits i.e., k
 );
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L0 ; // These wires are used to connect the outputs of each stage to the inputs of subsequent stages in the pipeline.
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L1 ; // L0 is output k bits of 1st stage, similarly L63 is output kbits of 64th stage
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L2 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L3 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L4 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L5 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L6 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L7 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L8 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L9 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L10 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L11 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L12 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L13 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L14 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L15 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L16 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L17 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L18 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L19 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L20 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L21 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L22 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L23 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L24 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L25 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L26 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L27 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L28 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L29 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L30 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L31 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L32 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L33 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L34 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L35 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L36 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L37 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L38 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L39 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L40 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L41 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L42 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L43 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L44 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L45 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L46 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L47 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L48 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L49 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L50 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L51 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L52 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L53 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L54 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L55 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L56 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L57 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L58 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L59 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L60 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L61 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L62 ; 
(* DONT_TOUCH= "TRUE" *)wire [3 :0] L63 ; 

 assign oTP = L63 ; 
 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage0( {4{itriger}},{4{itriger}}, iC[0], L0); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage1( { L0[3], L0[2], L0[0], L0[1]}, { L0[1], L0[0], L0[3], L0[2]}, iC[1],  L1); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage2( { L1[1], L1[2], L1[0], L1[3]}, { L1[0], L1[3], L1[2], L1[1]}, iC[2],  L2); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage3( { L2[1], L2[0], L2[3], L2[2]}, { L2[2], L2[3], L2[1], L2[0]}, iC[3],  L3); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage4( { L3[0], L3[3], L3[2], L3[1]}, { L3[1], L3[2], L3[3], L3[0]}, iC[4],  L4); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage5( { L4[3], L4[1], L4[2], L4[0]}, { L4[2], L4[0], L4[1], L4[3]}, iC[5],  L5); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage6( { L5[1], L5[3], L5[0], L5[2]}, { L5[2], L5[0], L5[1], L5[3]}, iC[6],  L6); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage7( { L6[0], L6[2], L6[1], L6[3]}, { L6[3], L6[0], L6[2], L6[1]}, iC[7],  L7); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage8( { L7[0], L7[2], L7[3], L7[1]}, { L7[1], L7[3], L7[0], L7[2]}, iC[8],  L8); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage9( { L8[0], L8[2], L8[3], L8[1]}, { L8[3], L8[1], L8[2], L8[0]}, iC[9],  L9); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage10( { L9[0], L9[3], L9[1], L9[2]}, { L9[2], L9[0], L9[3], L9[1]}, iC[10],  L10); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage11( { L10[1], L10[3], L10[0], L10[2]}, { L10[3], L10[2], L10[1], L10[0]}, iC[11],  L11); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage12( { L11[1], L11[3], L11[2], L11[0]}, { L11[0], L11[1], L11[3], L11[2]}, iC[12],  L12); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage13( { L12[1], L12[3], L12[2], L12[0]}, { L12[2], L12[0], L12[1], L12[3]}, iC[13],  L13); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage14( { L13[0], L13[2], L13[3], L13[1]}, { L13[3], L13[0], L13[1], L13[2]}, iC[14],  L14); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage15( { L14[3], L14[1], L14[2], L14[0]}, { L14[2], L14[0], L14[3], L14[1]}, iC[15],  L15); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage16( { L15[0], L15[1], L15[2], L15[3]}, { L15[3], L15[2], L15[0], L15[1]}, iC[16],  L16); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage17( { L16[0], L16[3], L16[1], L16[2]}, { L16[1], L16[2], L16[3], L16[0]}, iC[17],  L17); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage18( { L17[1], L17[0], L17[2], L17[3]}, { L17[2], L17[1], L17[3], L17[0]}, iC[18],  L18); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage19( { L18[2], L18[3], L18[1], L18[0]}, { L18[1], L18[2], L18[0], L18[3]}, iC[19],  L19); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage20( { L19[0], L19[3], L19[1], L19[2]}, { L19[2], L19[1], L19[3], L19[0]}, iC[20],  L20); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage21( { L20[2], L20[3], L20[0], L20[1]}, { L20[3], L20[2], L20[1], L20[0]}, iC[21],  L21); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage22( { L21[0], L21[1], L21[2], L21[3]}, { L21[3], L21[2], L21[0], L21[1]}, iC[22],  L22); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage23( { L22[3], L22[0], L22[2], L22[1]}, { L22[0], L22[1], L22[3], L22[2]}, iC[23],  L23); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage24( { L23[3], L23[1], L23[0], L23[2]}, { L23[1], L23[0], L23[2], L23[3]}, iC[24],  L24); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage25( { L24[3], L24[0], L24[2], L24[1]}, { L24[0], L24[2], L24[1], L24[3]}, iC[25],  L25); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage26( { L25[3], L25[0], L25[2], L25[1]}, { L25[1], L25[2], L25[0], L25[3]}, iC[26],  L26); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage27( { L26[0], L26[2], L26[3], L26[1]}, { L26[1], L26[0], L26[2], L26[3]}, iC[27],  L27); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage28( { L27[2], L27[3], L27[1], L27[0]}, { L27[0], L27[2], L27[3], L27[1]}, iC[28],  L28); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage29( { L28[0], L28[3], L28[1], L28[2]}, { L28[2], L28[1], L28[3], L28[0]}, iC[29],  L29); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage30( { L29[3], L29[1], L29[0], L29[2]}, { L29[0], L29[2], L29[1], L29[3]}, iC[30],  L30); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage31( { L30[1], L30[0], L30[2], L30[3]}, { L30[3], L30[2], L30[1], L30[0]}, iC[31],  L31); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage32( { L31[2], L31[3], L31[1], L31[0]}, { L31[1], L31[0], L31[2], L31[3]}, iC[32],  L32); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage33( { L32[3], L32[0], L32[1], L32[2]}, { L32[0], L32[2], L32[3], L32[1]}, iC[33],  L33); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage34( { L33[0], L33[3], L33[1], L33[2]}, { L33[3], L33[1], L33[2], L33[0]}, iC[34],  L34); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage35( { L34[1], L34[0], L34[3], L34[2]}, { L34[0], L34[3], L34[2], L34[1]}, iC[35],  L35); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage36( { L35[2], L35[1], L35[0], L35[3]}, { L35[0], L35[3], L35[1], L35[2]}, iC[36],  L36); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage37( { L36[1], L36[3], L36[2], L36[0]}, { L36[3], L36[2], L36[0], L36[1]}, iC[37],  L37); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage38( { L37[3], L37[2], L37[1], L37[0]}, { L37[2], L37[1], L37[0], L37[3]}, iC[38],  L38); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage39( { L38[2], L38[0], L38[1], L38[3]}, { L38[3], L38[1], L38[2], L38[0]}, iC[39],  L39); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage40( { L39[1], L39[3], L39[2], L39[0]}, { L39[2], L39[0], L39[3], L39[1]}, iC[40],  L40); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage41( { L40[2], L40[1], L40[3], L40[0]}, { L40[0], L40[2], L40[1], L40[3]}, iC[41],  L41); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage42( { L41[2], L41[3], L41[0], L41[1]}, { L41[3], L41[1], L41[2], L41[0]}, iC[42],  L42); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage43( { L42[1], L42[3], L42[2], L42[0]}, { L42[2], L42[1], L42[0], L42[3]}, iC[43],  L43); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage44( { L43[0], L43[1], L43[3], L43[2]}, { L43[3], L43[2], L43[0], L43[1]}, iC[44],  L44); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage45( { L44[1], L44[0], L44[3], L44[2]}, { L44[0], L44[1], L44[2], L44[3]}, iC[45],  L45); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage46( { L45[3], L45[2], L45[1], L45[0]}, { L45[1], L45[0], L45[2], L45[3]}, iC[46],  L46); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage47( { L46[3], L46[1], L46[2], L46[0]}, { L46[0], L46[2], L46[1], L46[3]}, iC[47],  L47); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage48( { L47[1], L47[0], L47[3], L47[2]}, { L47[0], L47[1], L47[2], L47[3]}, iC[48],  L48); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage49( { L48[1], L48[3], L48[0], L48[2]}, { L48[0], L48[2], L48[1], L48[3]}, iC[49],  L49); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage50( { L49[2], L49[0], L49[1], L49[3]}, { L49[3], L49[1], L49[0], L49[2]}, iC[50],  L50); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage51( { L50[3], L50[0], L50[2], L50[1]}, { L50[2], L50[1], L50[3], L50[0]}, iC[51],  L51); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage52( { L51[1], L51[0], L51[2], L51[3]}, { L51[3], L51[2], L51[0], L51[1]}, iC[52],  L52); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage53( { L52[2], L52[0], L52[1], L52[3]}, { L52[3], L52[1], L52[0], L52[2]}, iC[53],  L53); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage54( { L53[1], L53[3], L53[2], L53[0]}, { L53[3], L53[1], L53[0], L53[2]}, iC[54],  L54); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage55( { L54[0], L54[3], L54[2], L54[1]}, { L54[1], L54[0], L54[3], L54[2]}, iC[55],  L55); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage56( { L55[1], L55[2], L55[3], L55[0]}, { L55[0], L55[1], L55[2], L55[3]}, iC[56],  L56); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage57( { L56[0], L56[2], L56[1], L56[3]}, { L56[2], L56[0], L56[3], L56[1]}, iC[57],  L57); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage58( { L57[2], L57[0], L57[3], L57[1]}, { L57[1], L57[2], L57[0], L57[3]}, iC[58],  L58); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage59( { L58[1], L58[0], L58[3], L58[2]}, { L58[2], L58[3], L58[1], L58[0]}, iC[59],  L59); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage60( { L59[2], L59[3], L59[1], L59[0]}, { L59[3], L59[2], L59[0], L59[1]}, iC[60],  L60); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage61( { L60[3], L60[2], L60[1], L60[0]}, { L60[1], L60[0], L60[2], L60[3]}, iC[61],  L61); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage62( { L61[2], L61[1], L61[0], L61[3]}, { L61[1], L61[3], L61[2], L61[0]}, iC[62],  L62); 
(*KEEP_HIERARCHY = "TRUE"*) MUX2to1_group #(.DW(4)) stage63( { L62[2], L62[0], L62[3], L62[1]}, { L62[3], L62[1], L62[0], L62[2]}, iC[63],  L63); 

 endmodule 
